conectix             '��Xqemu  Wi2k                       ����~���MM�b^�&�m                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������conectix             '��Xqemu  Wi2k                       ����~���MM�b^�&�m                                                                                                                                                                                                                                                                                                                                                                                                                                            